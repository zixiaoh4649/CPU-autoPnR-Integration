/home/zixiaoh3/ece425/pnr_provide/stdcells.lef
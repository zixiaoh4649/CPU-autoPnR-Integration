/home/zixiaoh3/ece425.work/pnr_provide/regfile.lef
/home/zixiaoh3/Desktop/backup/pnr/pnr_cpu1_success/pnr_provide/stdcells.lef